module tb_hack_top();

// Inputs
reg clk;
reg reset;

// Instantiate the hack_top module
hack_top dut (
.clk(clk),
.reset(reset)
);

logic [16384 -1 :0][15:0] mem;
// Clock generation
always #5 clk = ~clk;


always @(*)begin
/* using instance of mem to reflect a memory

msb = 7
lsb = 0

# Open the file in write mode
file = open('text_for_testbench_top_hack.txt', 'w')

# Loop through the ranges and write each value of s to the file
for a in range(4):
    for b in range(8):
        for c in range(8):
            for d in range(8):
                s = f"mem[{msb}:{lsb}] = dut.ram16k_inst.genblk1[{a}].ram4k_inst.genblk1[{b}].ram512_inst.genblk1[{c}].ram64_inst.genblk1[{d}].ram8_inst.mem;"
                file.write(s + "\n")

                # Update msb and lsb
                msb += 8
                lsb += 8

# Close the file
file.close()

*/
 mem[7:0]  =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[15:8] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[23:16] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[31:24] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[39:32] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[47:40] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[55:48] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[63:56] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[71:64] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[79:72] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[87:80] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[95:88] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[103:96] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[111:104] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[119:112] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[127:120] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[135:128] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[143:136] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[151:144] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[159:152] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[167:160] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[175:168] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[183:176] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[191:184] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[199:192] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[207:200] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[215:208] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[223:216] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[231:224] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[239:232] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[247:240] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[255:248] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[263:256] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[271:264] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[279:272] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[287:280] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[295:288] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[303:296] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[311:304] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[319:312] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[327:320] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[335:328] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[343:336] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[351:344] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[359:352] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[367:360] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[375:368] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[383:376] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[391:384] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[399:392] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[407:400] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[415:408] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[423:416] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[431:424] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[439:432] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[447:440] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[455:448] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[463:456] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[471:464] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[479:472] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[487:480] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[495:488] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[503:496] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[511:504] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[519:512] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[527:520] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[535:528] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[543:536] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[551:544] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[559:552] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[567:560] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[575:568] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[583:576] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[591:584] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[599:592] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[607:600] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[615:608] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[623:616] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[631:624] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[639:632] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[647:640] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[655:648] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[663:656] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[671:664] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[679:672] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[687:680] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[695:688] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[703:696] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[711:704] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[719:712] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[727:720] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[735:728] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[743:736] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[751:744] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[759:752] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[767:760] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[775:768] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[783:776] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[791:784] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[799:792] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[807:800] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[815:808] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[823:816] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[831:824] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[839:832] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[847:840] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[855:848] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[863:856] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[871:864] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[879:872] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[887:880] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[895:888] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[903:896] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[911:904] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[919:912] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[927:920] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[935:928] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[943:936] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[951:944] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[959:952] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[967:960] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[975:968] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[983:976] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[991:984] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[999:992] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[1007:1000] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[1015:1008] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[1023:1016] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[1031:1024] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[1039:1032] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[1047:1040] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[1055:1048] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[1063:1056] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[1071:1064] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[1079:1072] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[1087:1080] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[1095:1088] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[1103:1096] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[1111:1104] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[1119:1112] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[1127:1120] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[1135:1128] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[1143:1136] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[1151:1144] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[1159:1152] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[1167:1160] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[1175:1168] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[1183:1176] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[1191:1184] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[1199:1192] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[1207:1200] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[1215:1208] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[1223:1216] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[1231:1224] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[1239:1232] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[1247:1240] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[1255:1248] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[1263:1256] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[1271:1264] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[1279:1272] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[1287:1280] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[1295:1288] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[1303:1296] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[1311:1304] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[1319:1312] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[1327:1320] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[1335:1328] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[1343:1336] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[1351:1344] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[1359:1352] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[1367:1360] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[1375:1368] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[1383:1376] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[1391:1384] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[1399:1392] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[1407:1400] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[1415:1408] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[1423:1416] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[1431:1424] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[1439:1432] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[1447:1440] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[1455:1448] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[1463:1456] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[1471:1464] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[1479:1472] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[1487:1480] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[1495:1488] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[1503:1496] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[1511:1504] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[1519:1512] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[1527:1520] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[1535:1528] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[1543:1536] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[1551:1544] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[1559:1552] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[1567:1560] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[1575:1568] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[1583:1576] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[1591:1584] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[1599:1592] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[1607:1600] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[1615:1608] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[1623:1616] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[1631:1624] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[1639:1632] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[1647:1640] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[1655:1648] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[1663:1656] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[1671:1664] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[1679:1672] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[1687:1680] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[1695:1688] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[1703:1696] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[1711:1704] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[1719:1712] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[1727:1720] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[1735:1728] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[1743:1736] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[1751:1744] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[1759:1752] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[1767:1760] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[1775:1768] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[1783:1776] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[1791:1784] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[1799:1792] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[1807:1800] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[1815:1808] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[1823:1816] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[1831:1824] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[1839:1832] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[1847:1840] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[1855:1848] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[1863:1856] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[1871:1864] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[1879:1872] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[1887:1880] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[1895:1888] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[1903:1896] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[1911:1904] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[1919:1912] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[1927:1920] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[1935:1928] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[1943:1936] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[1951:1944] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[1959:1952] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[1967:1960] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[1975:1968] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[1983:1976] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[1991:1984] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[1999:1992] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[2007:2000] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[2015:2008] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[2023:2016] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[2031:2024] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[2039:2032] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[2047:2040] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[2055:2048] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[2063:2056] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[2071:2064] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[2079:2072] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[2087:2080] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[2095:2088] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[2103:2096] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[2111:2104] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[2119:2112] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[2127:2120] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[2135:2128] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[2143:2136] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[2151:2144] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[2159:2152] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[2167:2160] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[2175:2168] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[2183:2176] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[2191:2184] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[2199:2192] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[2207:2200] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[2215:2208] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[2223:2216] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[2231:2224] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[2239:2232] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[2247:2240] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[2255:2248] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[2263:2256] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[2271:2264] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[2279:2272] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[2287:2280] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[2295:2288] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[2303:2296] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[2311:2304] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[2319:2312] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[2327:2320] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[2335:2328] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[2343:2336] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[2351:2344] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[2359:2352] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[2367:2360] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[2375:2368] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[2383:2376] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[2391:2384] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[2399:2392] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[2407:2400] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[2415:2408] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[2423:2416] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[2431:2424] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[2439:2432] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[2447:2440] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[2455:2448] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[2463:2456] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[2471:2464] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[2479:2472] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[2487:2480] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[2495:2488] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[2503:2496] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[2511:2504] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[2519:2512] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[2527:2520] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[2535:2528] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[2543:2536] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[2551:2544] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[2559:2552] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[2567:2560] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[2575:2568] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[2583:2576] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[2591:2584] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[2599:2592] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[2607:2600] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[2615:2608] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[2623:2616] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[2631:2624] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[2639:2632] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[2647:2640] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[2655:2648] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[2663:2656] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[2671:2664] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[2679:2672] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[2687:2680] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[2695:2688] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[2703:2696] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[2711:2704] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[2719:2712] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[2727:2720] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[2735:2728] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[2743:2736] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[2751:2744] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[2759:2752] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[2767:2760] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[2775:2768] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[2783:2776] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[2791:2784] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[2799:2792] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[2807:2800] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[2815:2808] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[2823:2816] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[2831:2824] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[2839:2832] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[2847:2840] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[2855:2848] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[2863:2856] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[2871:2864] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[2879:2872] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[2887:2880] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[2895:2888] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[2903:2896] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[2911:2904] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[2919:2912] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[2927:2920] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[2935:2928] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[2943:2936] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[2951:2944] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[2959:2952] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[2967:2960] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[2975:2968] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[2983:2976] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[2991:2984] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[2999:2992] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[3007:3000] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[3015:3008] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[3023:3016] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[3031:3024] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[3039:3032] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[3047:3040] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[3055:3048] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[3063:3056] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[3071:3064] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[3079:3072] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[3087:3080] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[3095:3088] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[3103:3096] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[3111:3104] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[3119:3112] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[3127:3120] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[3135:3128] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[3143:3136] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[3151:3144] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[3159:3152] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[3167:3160] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[3175:3168] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[3183:3176] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[3191:3184] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[3199:3192] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[3207:3200] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[3215:3208] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[3223:3216] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[3231:3224] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[3239:3232] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[3247:3240] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[3255:3248] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[3263:3256] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[3271:3264] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[3279:3272] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[3287:3280] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[3295:3288] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[3303:3296] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[3311:3304] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[3319:3312] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[3327:3320] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[3335:3328] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[3343:3336] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[3351:3344] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[3359:3352] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[3367:3360] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[3375:3368] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[3383:3376] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[3391:3384] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[3399:3392] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[3407:3400] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[3415:3408] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[3423:3416] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[3431:3424] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[3439:3432] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[3447:3440] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[3455:3448] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[3463:3456] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[3471:3464] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[3479:3472] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[3487:3480] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[3495:3488] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[3503:3496] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[3511:3504] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[3519:3512] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[3527:3520] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[3535:3528] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[3543:3536] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[3551:3544] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[3559:3552] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[3567:3560] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[3575:3568] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[3583:3576] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[3591:3584] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[3599:3592] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[3607:3600] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[3615:3608] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[3623:3616] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[3631:3624] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[3639:3632] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[3647:3640] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[3655:3648] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[3663:3656] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[3671:3664] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[3679:3672] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[3687:3680] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[3695:3688] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[3703:3696] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[3711:3704] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[3719:3712] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[3727:3720] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[3735:3728] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[3743:3736] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[3751:3744] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[3759:3752] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[3767:3760] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[3775:3768] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[3783:3776] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[3791:3784] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[3799:3792] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[3807:3800] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[3815:3808] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[3823:3816] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[3831:3824] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[3839:3832] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[3847:3840] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[3855:3848] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[3863:3856] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[3871:3864] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[3879:3872] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[3887:3880] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[3895:3888] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[3903:3896] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[3911:3904] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[3919:3912] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[3927:3920] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[3935:3928] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[3943:3936] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[3951:3944] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[3959:3952] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[3967:3960] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[3975:3968] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[3983:3976] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[3991:3984] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[3999:3992] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[4007:4000] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[4015:4008] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[4023:4016] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[4031:4024] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[4039:4032] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[4047:4040] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[4055:4048] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[4063:4056] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[4071:4064] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[4079:4072] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[4087:4080] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[4095:4088] =dut.ram16k_inst.genblk1[0].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[4103:4096] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[4111:4104] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[4119:4112] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[4127:4120] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[4135:4128] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[4143:4136] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[4151:4144] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[4159:4152] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[4167:4160] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[4175:4168] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[4183:4176] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[4191:4184] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[4199:4192] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[4207:4200] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[4215:4208] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[4223:4216] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[4231:4224] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[4239:4232] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[4247:4240] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[4255:4248] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[4263:4256] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[4271:4264] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[4279:4272] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[4287:4280] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[4295:4288] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[4303:4296] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[4311:4304] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[4319:4312] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[4327:4320] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[4335:4328] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[4343:4336] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[4351:4344] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[4359:4352] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[4367:4360] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[4375:4368] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[4383:4376] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[4391:4384] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[4399:4392] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[4407:4400] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[4415:4408] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[4423:4416] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[4431:4424] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[4439:4432] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[4447:4440] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[4455:4448] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[4463:4456] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[4471:4464] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[4479:4472] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[4487:4480] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[4495:4488] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[4503:4496] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[4511:4504] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[4519:4512] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[4527:4520] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[4535:4528] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[4543:4536] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[4551:4544] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[4559:4552] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[4567:4560] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[4575:4568] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[4583:4576] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[4591:4584] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[4599:4592] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[4607:4600] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[4615:4608] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[4623:4616] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[4631:4624] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[4639:4632] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[4647:4640] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[4655:4648] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[4663:4656] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[4671:4664] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[4679:4672] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[4687:4680] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[4695:4688] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[4703:4696] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[4711:4704] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[4719:4712] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[4727:4720] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[4735:4728] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[4743:4736] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[4751:4744] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[4759:4752] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[4767:4760] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[4775:4768] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[4783:4776] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[4791:4784] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[4799:4792] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[4807:4800] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[4815:4808] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[4823:4816] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[4831:4824] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[4839:4832] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[4847:4840] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[4855:4848] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[4863:4856] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[4871:4864] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[4879:4872] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[4887:4880] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[4895:4888] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[4903:4896] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[4911:4904] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[4919:4912] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[4927:4920] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[4935:4928] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[4943:4936] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[4951:4944] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[4959:4952] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[4967:4960] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[4975:4968] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[4983:4976] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[4991:4984] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[4999:4992] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[5007:5000] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[5015:5008] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[5023:5016] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[5031:5024] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[5039:5032] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[5047:5040] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[5055:5048] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[5063:5056] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[5071:5064] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[5079:5072] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[5087:5080] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[5095:5088] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[5103:5096] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[5111:5104] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[5119:5112] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[5127:5120] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[5135:5128] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[5143:5136] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[5151:5144] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[5159:5152] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[5167:5160] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[5175:5168] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[5183:5176] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[5191:5184] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[5199:5192] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[5207:5200] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[5215:5208] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[5223:5216] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[5231:5224] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[5239:5232] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[5247:5240] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[5255:5248] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[5263:5256] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[5271:5264] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[5279:5272] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[5287:5280] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[5295:5288] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[5303:5296] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[5311:5304] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[5319:5312] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[5327:5320] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[5335:5328] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[5343:5336] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[5351:5344] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[5359:5352] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[5367:5360] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[5375:5368] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[5383:5376] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[5391:5384] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[5399:5392] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[5407:5400] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[5415:5408] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[5423:5416] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[5431:5424] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[5439:5432] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[5447:5440] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[5455:5448] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[5463:5456] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[5471:5464] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[5479:5472] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[5487:5480] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[5495:5488] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[5503:5496] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[5511:5504] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[5519:5512] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[5527:5520] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[5535:5528] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[5543:5536] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[5551:5544] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[5559:5552] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[5567:5560] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[5575:5568] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[5583:5576] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[5591:5584] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[5599:5592] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[5607:5600] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[5615:5608] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[5623:5616] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[5631:5624] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[5639:5632] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[5647:5640] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[5655:5648] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[5663:5656] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[5671:5664] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[5679:5672] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[5687:5680] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[5695:5688] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[5703:5696] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[5711:5704] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[5719:5712] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[5727:5720] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[5735:5728] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[5743:5736] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[5751:5744] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[5759:5752] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[5767:5760] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[5775:5768] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[5783:5776] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[5791:5784] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[5799:5792] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[5807:5800] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[5815:5808] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[5823:5816] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[5831:5824] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[5839:5832] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[5847:5840] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[5855:5848] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[5863:5856] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[5871:5864] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[5879:5872] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[5887:5880] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[5895:5888] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[5903:5896] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[5911:5904] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[5919:5912] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[5927:5920] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[5935:5928] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[5943:5936] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[5951:5944] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[5959:5952] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[5967:5960] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[5975:5968] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[5983:5976] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[5991:5984] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[5999:5992] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[6007:6000] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[6015:6008] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[6023:6016] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[6031:6024] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[6039:6032] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[6047:6040] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[6055:6048] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[6063:6056] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[6071:6064] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[6079:6072] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[6087:6080] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[6095:6088] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[6103:6096] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[6111:6104] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[6119:6112] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[6127:6120] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[6135:6128] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[6143:6136] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[6151:6144] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[6159:6152] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[6167:6160] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[6175:6168] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[6183:6176] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[6191:6184] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[6199:6192] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[6207:6200] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[6215:6208] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[6223:6216] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[6231:6224] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[6239:6232] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[6247:6240] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[6255:6248] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[6263:6256] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[6271:6264] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[6279:6272] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[6287:6280] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[6295:6288] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[6303:6296] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[6311:6304] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[6319:6312] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[6327:6320] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[6335:6328] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[6343:6336] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[6351:6344] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[6359:6352] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[6367:6360] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[6375:6368] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[6383:6376] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[6391:6384] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[6399:6392] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[6407:6400] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[6415:6408] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[6423:6416] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[6431:6424] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[6439:6432] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[6447:6440] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[6455:6448] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[6463:6456] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[6471:6464] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[6479:6472] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[6487:6480] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[6495:6488] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[6503:6496] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[6511:6504] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[6519:6512] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[6527:6520] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[6535:6528] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[6543:6536] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[6551:6544] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[6559:6552] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[6567:6560] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[6575:6568] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[6583:6576] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[6591:6584] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[6599:6592] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[6607:6600] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[6615:6608] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[6623:6616] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[6631:6624] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[6639:6632] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[6647:6640] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[6655:6648] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[6663:6656] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[6671:6664] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[6679:6672] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[6687:6680] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[6695:6688] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[6703:6696] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[6711:6704] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[6719:6712] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[6727:6720] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[6735:6728] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[6743:6736] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[6751:6744] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[6759:6752] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[6767:6760] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[6775:6768] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[6783:6776] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[6791:6784] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[6799:6792] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[6807:6800] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[6815:6808] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[6823:6816] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[6831:6824] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[6839:6832] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[6847:6840] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[6855:6848] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[6863:6856] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[6871:6864] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[6879:6872] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[6887:6880] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[6895:6888] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[6903:6896] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[6911:6904] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[6919:6912] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[6927:6920] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[6935:6928] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[6943:6936] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[6951:6944] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[6959:6952] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[6967:6960] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[6975:6968] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[6983:6976] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[6991:6984] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[6999:6992] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[7007:7000] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[7015:7008] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[7023:7016] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[7031:7024] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[7039:7032] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[7047:7040] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[7055:7048] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[7063:7056] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[7071:7064] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[7079:7072] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[7087:7080] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[7095:7088] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[7103:7096] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[7111:7104] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[7119:7112] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[7127:7120] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[7135:7128] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[7143:7136] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[7151:7144] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[7159:7152] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[7167:7160] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[7175:7168] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[7183:7176] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[7191:7184] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[7199:7192] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[7207:7200] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[7215:7208] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[7223:7216] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[7231:7224] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[7239:7232] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[7247:7240] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[7255:7248] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[7263:7256] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[7271:7264] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[7279:7272] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[7287:7280] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[7295:7288] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[7303:7296] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[7311:7304] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[7319:7312] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[7327:7320] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[7335:7328] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[7343:7336] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[7351:7344] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[7359:7352] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[7367:7360] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[7375:7368] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[7383:7376] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[7391:7384] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[7399:7392] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[7407:7400] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[7415:7408] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[7423:7416] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[7431:7424] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[7439:7432] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[7447:7440] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[7455:7448] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[7463:7456] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[7471:7464] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[7479:7472] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[7487:7480] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[7495:7488] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[7503:7496] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[7511:7504] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[7519:7512] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[7527:7520] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[7535:7528] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[7543:7536] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[7551:7544] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[7559:7552] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[7567:7560] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[7575:7568] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[7583:7576] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[7591:7584] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[7599:7592] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[7607:7600] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[7615:7608] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[7623:7616] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[7631:7624] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[7639:7632] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[7647:7640] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[7655:7648] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[7663:7656] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[7671:7664] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[7679:7672] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[7687:7680] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[7695:7688] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[7703:7696] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[7711:7704] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[7719:7712] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[7727:7720] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[7735:7728] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[7743:7736] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[7751:7744] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[7759:7752] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[7767:7760] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[7775:7768] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[7783:7776] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[7791:7784] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[7799:7792] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[7807:7800] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[7815:7808] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[7823:7816] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[7831:7824] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[7839:7832] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[7847:7840] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[7855:7848] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[7863:7856] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[7871:7864] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[7879:7872] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[7887:7880] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[7895:7888] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[7903:7896] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[7911:7904] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[7919:7912] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[7927:7920] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[7935:7928] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[7943:7936] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[7951:7944] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[7959:7952] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[7967:7960] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[7975:7968] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[7983:7976] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[7991:7984] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[7999:7992] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[8007:8000] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[8015:8008] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[8023:8016] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[8031:8024] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[8039:8032] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[8047:8040] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[8055:8048] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[8063:8056] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[8071:8064] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[8079:8072] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[8087:8080] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[8095:8088] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[8103:8096] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[8111:8104] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[8119:8112] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[8127:8120] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[8135:8128] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[8143:8136] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[8151:8144] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[8159:8152] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[8167:8160] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[8175:8168] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[8183:8176] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[8191:8184] =dut.ram16k_inst.genblk1[1].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[8199:8192] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[8207:8200] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[8215:8208] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[8223:8216] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[8231:8224] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[8239:8232] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[8247:8240] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[8255:8248] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[8263:8256] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[8271:8264] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[8279:8272] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[8287:8280] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[8295:8288] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[8303:8296] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[8311:8304] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[8319:8312] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[8327:8320] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[8335:8328] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[8343:8336] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[8351:8344] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[8359:8352] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[8367:8360] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[8375:8368] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[8383:8376] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[8391:8384] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[8399:8392] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[8407:8400] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[8415:8408] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[8423:8416] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[8431:8424] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[8439:8432] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[8447:8440] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[8455:8448] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[8463:8456] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[8471:8464] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[8479:8472] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[8487:8480] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[8495:8488] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[8503:8496] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[8511:8504] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[8519:8512] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[8527:8520] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[8535:8528] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[8543:8536] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[8551:8544] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[8559:8552] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[8567:8560] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[8575:8568] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[8583:8576] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[8591:8584] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[8599:8592] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[8607:8600] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[8615:8608] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[8623:8616] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[8631:8624] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[8639:8632] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[8647:8640] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[8655:8648] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[8663:8656] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[8671:8664] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[8679:8672] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[8687:8680] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[8695:8688] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[8703:8696] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[8711:8704] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[8719:8712] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[8727:8720] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[8735:8728] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[8743:8736] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[8751:8744] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[8759:8752] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[8767:8760] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[8775:8768] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[8783:8776] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[8791:8784] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[8799:8792] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[8807:8800] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[8815:8808] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[8823:8816] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[8831:8824] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[8839:8832] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[8847:8840] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[8855:8848] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[8863:8856] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[8871:8864] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[8879:8872] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[8887:8880] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[8895:8888] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[8903:8896] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[8911:8904] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[8919:8912] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[8927:8920] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[8935:8928] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[8943:8936] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[8951:8944] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[8959:8952] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[8967:8960] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[8975:8968] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[8983:8976] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[8991:8984] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[8999:8992] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[9007:9000] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[9015:9008] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[9023:9016] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[9031:9024] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[9039:9032] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[9047:9040] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[9055:9048] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[9063:9056] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[9071:9064] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[9079:9072] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[9087:9080] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[9095:9088] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[9103:9096] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[9111:9104] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[9119:9112] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[9127:9120] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[9135:9128] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[9143:9136] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[9151:9144] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[9159:9152] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[9167:9160] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[9175:9168] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[9183:9176] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[9191:9184] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[9199:9192] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[9207:9200] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[9215:9208] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[9223:9216] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[9231:9224] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[9239:9232] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[9247:9240] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[9255:9248] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[9263:9256] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[9271:9264] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[9279:9272] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[9287:9280] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[9295:9288] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[9303:9296] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[9311:9304] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[9319:9312] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[9327:9320] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[9335:9328] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[9343:9336] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[9351:9344] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[9359:9352] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[9367:9360] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[9375:9368] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[9383:9376] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[9391:9384] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[9399:9392] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[9407:9400] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[9415:9408] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[9423:9416] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[9431:9424] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[9439:9432] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[9447:9440] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[9455:9448] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[9463:9456] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[9471:9464] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[9479:9472] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[9487:9480] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[9495:9488] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[9503:9496] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[9511:9504] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[9519:9512] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[9527:9520] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[9535:9528] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[9543:9536] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[9551:9544] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[9559:9552] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[9567:9560] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[9575:9568] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[9583:9576] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[9591:9584] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[9599:9592] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[9607:9600] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[9615:9608] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[9623:9616] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[9631:9624] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[9639:9632] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[9647:9640] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[9655:9648] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[9663:9656] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[9671:9664] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[9679:9672] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[9687:9680] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[9695:9688] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[9703:9696] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[9711:9704] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[9719:9712] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[9727:9720] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[9735:9728] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[9743:9736] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[9751:9744] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[9759:9752] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[9767:9760] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[9775:9768] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[9783:9776] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[9791:9784] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[9799:9792] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[9807:9800] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[9815:9808] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[9823:9816] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[9831:9824] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[9839:9832] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[9847:9840] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[9855:9848] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[9863:9856] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[9871:9864] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[9879:9872] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[9887:9880] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[9895:9888] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[9903:9896] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[9911:9904] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[9919:9912] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[9927:9920] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[9935:9928] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[9943:9936] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[9951:9944] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[9959:9952] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[9967:9960] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[9975:9968] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[9983:9976] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[9991:9984] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[9999:9992] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[10007:10000] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[10015:10008] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[10023:10016] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[10031:10024] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[10039:10032] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[10047:10040] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[10055:10048] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[10063:10056] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[10071:10064] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[10079:10072] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[10087:10080] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[10095:10088] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[10103:10096] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[10111:10104] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[10119:10112] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[10127:10120] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[10135:10128] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[10143:10136] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[10151:10144] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[10159:10152] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[10167:10160] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[10175:10168] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[10183:10176] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[10191:10184] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[10199:10192] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[10207:10200] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[10215:10208] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[10223:10216] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[10231:10224] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[10239:10232] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[10247:10240] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[10255:10248] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[10263:10256] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[10271:10264] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[10279:10272] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[10287:10280] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[10295:10288] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[10303:10296] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[10311:10304] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[10319:10312] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[10327:10320] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[10335:10328] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[10343:10336] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[10351:10344] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[10359:10352] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[10367:10360] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[10375:10368] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[10383:10376] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[10391:10384] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[10399:10392] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[10407:10400] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[10415:10408] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[10423:10416] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[10431:10424] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[10439:10432] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[10447:10440] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[10455:10448] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[10463:10456] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[10471:10464] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[10479:10472] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[10487:10480] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[10495:10488] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[10503:10496] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[10511:10504] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[10519:10512] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[10527:10520] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[10535:10528] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[10543:10536] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[10551:10544] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[10559:10552] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[10567:10560] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[10575:10568] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[10583:10576] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[10591:10584] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[10599:10592] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[10607:10600] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[10615:10608] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[10623:10616] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[10631:10624] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[10639:10632] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[10647:10640] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[10655:10648] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[10663:10656] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[10671:10664] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[10679:10672] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[10687:10680] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[10695:10688] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[10703:10696] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[10711:10704] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[10719:10712] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[10727:10720] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[10735:10728] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[10743:10736] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[10751:10744] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[10759:10752] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[10767:10760] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[10775:10768] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[10783:10776] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[10791:10784] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[10799:10792] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[10807:10800] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[10815:10808] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[10823:10816] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[10831:10824] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[10839:10832] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[10847:10840] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[10855:10848] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[10863:10856] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[10871:10864] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[10879:10872] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[10887:10880] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[10895:10888] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[10903:10896] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[10911:10904] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[10919:10912] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[10927:10920] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[10935:10928] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[10943:10936] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[10951:10944] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[10959:10952] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[10967:10960] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[10975:10968] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[10983:10976] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[10991:10984] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[10999:10992] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[11007:11000] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[11015:11008] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[11023:11016] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[11031:11024] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[11039:11032] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[11047:11040] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[11055:11048] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[11063:11056] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[11071:11064] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[11079:11072] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[11087:11080] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[11095:11088] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[11103:11096] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[11111:11104] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[11119:11112] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[11127:11120] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[11135:11128] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[11143:11136] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[11151:11144] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[11159:11152] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[11167:11160] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[11175:11168] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[11183:11176] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[11191:11184] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[11199:11192] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[11207:11200] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[11215:11208] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[11223:11216] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[11231:11224] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[11239:11232] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[11247:11240] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[11255:11248] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[11263:11256] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[11271:11264] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[11279:11272] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[11287:11280] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[11295:11288] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[11303:11296] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[11311:11304] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[11319:11312] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[11327:11320] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[11335:11328] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[11343:11336] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[11351:11344] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[11359:11352] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[11367:11360] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[11375:11368] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[11383:11376] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[11391:11384] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[11399:11392] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[11407:11400] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[11415:11408] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[11423:11416] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[11431:11424] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[11439:11432] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[11447:11440] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[11455:11448] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[11463:11456] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[11471:11464] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[11479:11472] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[11487:11480] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[11495:11488] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[11503:11496] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[11511:11504] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[11519:11512] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[11527:11520] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[11535:11528] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[11543:11536] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[11551:11544] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[11559:11552] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[11567:11560] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[11575:11568] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[11583:11576] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[11591:11584] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[11599:11592] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[11607:11600] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[11615:11608] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[11623:11616] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[11631:11624] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[11639:11632] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[11647:11640] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[11655:11648] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[11663:11656] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[11671:11664] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[11679:11672] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[11687:11680] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[11695:11688] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[11703:11696] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[11711:11704] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[11719:11712] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[11727:11720] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[11735:11728] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[11743:11736] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[11751:11744] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[11759:11752] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[11767:11760] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[11775:11768] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[11783:11776] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[11791:11784] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[11799:11792] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[11807:11800] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[11815:11808] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[11823:11816] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[11831:11824] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[11839:11832] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[11847:11840] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[11855:11848] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[11863:11856] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[11871:11864] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[11879:11872] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[11887:11880] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[11895:11888] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[11903:11896] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[11911:11904] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[11919:11912] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[11927:11920] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[11935:11928] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[11943:11936] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[11951:11944] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[11959:11952] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[11967:11960] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[11975:11968] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[11983:11976] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[11991:11984] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[11999:11992] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[12007:12000] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[12015:12008] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[12023:12016] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[12031:12024] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[12039:12032] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[12047:12040] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[12055:12048] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[12063:12056] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[12071:12064] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[12079:12072] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[12087:12080] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[12095:12088] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[12103:12096] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[12111:12104] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[12119:12112] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[12127:12120] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[12135:12128] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[12143:12136] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[12151:12144] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[12159:12152] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[12167:12160] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[12175:12168] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[12183:12176] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[12191:12184] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[12199:12192] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[12207:12200] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[12215:12208] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[12223:12216] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[12231:12224] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[12239:12232] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[12247:12240] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[12255:12248] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[12263:12256] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[12271:12264] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[12279:12272] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[12287:12280] =dut.ram16k_inst.genblk1[2].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[12295:12288] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[12303:12296] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[12311:12304] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[12319:12312] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[12327:12320] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[12335:12328] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[12343:12336] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[12351:12344] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[12359:12352] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[12367:12360] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[12375:12368] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[12383:12376] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[12391:12384] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[12399:12392] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[12407:12400] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[12415:12408] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[12423:12416] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[12431:12424] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[12439:12432] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[12447:12440] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[12455:12448] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[12463:12456] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[12471:12464] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[12479:12472] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[12487:12480] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[12495:12488] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[12503:12496] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[12511:12504] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[12519:12512] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[12527:12520] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[12535:12528] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[12543:12536] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[12551:12544] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[12559:12552] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[12567:12560] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[12575:12568] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[12583:12576] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[12591:12584] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[12599:12592] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[12607:12600] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[12615:12608] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[12623:12616] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[12631:12624] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[12639:12632] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[12647:12640] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[12655:12648] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[12663:12656] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[12671:12664] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[12679:12672] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[12687:12680] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[12695:12688] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[12703:12696] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[12711:12704] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[12719:12712] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[12727:12720] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[12735:12728] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[12743:12736] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[12751:12744] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[12759:12752] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[12767:12760] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[12775:12768] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[12783:12776] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[12791:12784] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[12799:12792] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[0].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[12807:12800] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[12815:12808] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[12823:12816] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[12831:12824] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[12839:12832] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[12847:12840] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[12855:12848] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[12863:12856] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[12871:12864] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[12879:12872] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[12887:12880] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[12895:12888] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[12903:12896] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[12911:12904] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[12919:12912] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[12927:12920] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[12935:12928] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[12943:12936] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[12951:12944] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[12959:12952] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[12967:12960] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[12975:12968] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[12983:12976] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[12991:12984] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[12999:12992] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[13007:13000] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[13015:13008] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[13023:13016] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[13031:13024] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[13039:13032] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[13047:13040] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[13055:13048] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[13063:13056] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[13071:13064] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[13079:13072] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[13087:13080] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[13095:13088] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[13103:13096] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[13111:13104] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[13119:13112] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[13127:13120] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[13135:13128] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[13143:13136] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[13151:13144] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[13159:13152] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[13167:13160] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[13175:13168] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[13183:13176] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[13191:13184] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[13199:13192] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[13207:13200] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[13215:13208] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[13223:13216] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[13231:13224] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[13239:13232] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[13247:13240] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[13255:13248] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[13263:13256] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[13271:13264] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[13279:13272] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[13287:13280] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[13295:13288] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[13303:13296] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[13311:13304] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[1].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[13319:13312] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[13327:13320] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[13335:13328] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[13343:13336] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[13351:13344] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[13359:13352] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[13367:13360] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[13375:13368] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[13383:13376] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[13391:13384] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[13399:13392] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[13407:13400] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[13415:13408] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[13423:13416] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[13431:13424] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[13439:13432] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[13447:13440] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[13455:13448] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[13463:13456] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[13471:13464] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[13479:13472] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[13487:13480] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[13495:13488] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[13503:13496] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[13511:13504] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[13519:13512] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[13527:13520] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[13535:13528] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[13543:13536] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[13551:13544] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[13559:13552] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[13567:13560] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[13575:13568] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[13583:13576] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[13591:13584] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[13599:13592] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[13607:13600] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[13615:13608] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[13623:13616] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[13631:13624] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[13639:13632] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[13647:13640] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[13655:13648] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[13663:13656] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[13671:13664] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[13679:13672] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[13687:13680] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[13695:13688] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[13703:13696] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[13711:13704] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[13719:13712] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[13727:13720] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[13735:13728] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[13743:13736] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[13751:13744] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[13759:13752] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[13767:13760] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[13775:13768] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[13783:13776] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[13791:13784] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[13799:13792] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[13807:13800] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[13815:13808] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[13823:13816] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[2].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[13831:13824] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[13839:13832] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[13847:13840] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[13855:13848] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[13863:13856] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[13871:13864] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[13879:13872] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[13887:13880] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[13895:13888] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[13903:13896] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[13911:13904] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[13919:13912] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[13927:13920] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[13935:13928] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[13943:13936] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[13951:13944] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[13959:13952] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[13967:13960] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[13975:13968] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[13983:13976] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[13991:13984] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[13999:13992] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[14007:14000] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[14015:14008] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[14023:14016] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[14031:14024] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[14039:14032] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[14047:14040] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[14055:14048] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[14063:14056] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[14071:14064] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[14079:14072] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[14087:14080] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[14095:14088] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[14103:14096] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[14111:14104] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[14119:14112] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[14127:14120] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[14135:14128] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[14143:14136] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[14151:14144] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[14159:14152] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[14167:14160] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[14175:14168] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[14183:14176] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[14191:14184] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[14199:14192] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[14207:14200] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[14215:14208] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[14223:14216] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[14231:14224] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[14239:14232] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[14247:14240] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[14255:14248] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[14263:14256] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[14271:14264] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[14279:14272] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[14287:14280] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[14295:14288] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[14303:14296] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[14311:14304] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[14319:14312] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[14327:14320] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[14335:14328] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[3].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[14343:14336] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[14351:14344] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[14359:14352] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[14367:14360] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[14375:14368] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[14383:14376] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[14391:14384] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[14399:14392] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[14407:14400] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[14415:14408] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[14423:14416] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[14431:14424] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[14439:14432] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[14447:14440] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[14455:14448] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[14463:14456] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[14471:14464] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[14479:14472] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[14487:14480] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[14495:14488] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[14503:14496] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[14511:14504] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[14519:14512] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[14527:14520] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[14535:14528] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[14543:14536] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[14551:14544] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[14559:14552] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[14567:14560] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[14575:14568] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[14583:14576] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[14591:14584] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[14599:14592] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[14607:14600] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[14615:14608] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[14623:14616] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[14631:14624] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[14639:14632] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[14647:14640] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[14655:14648] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[14663:14656] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[14671:14664] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[14679:14672] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[14687:14680] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[14695:14688] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[14703:14696] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[14711:14704] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[14719:14712] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[14727:14720] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[14735:14728] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[14743:14736] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[14751:14744] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[14759:14752] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[14767:14760] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[14775:14768] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[14783:14776] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[14791:14784] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[14799:14792] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[14807:14800] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[14815:14808] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[14823:14816] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[14831:14824] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[14839:14832] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[14847:14840] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[4].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[14855:14848] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[14863:14856] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[14871:14864] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[14879:14872] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[14887:14880] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[14895:14888] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[14903:14896] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[14911:14904] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[14919:14912] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[14927:14920] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[14935:14928] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[14943:14936] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[14951:14944] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[14959:14952] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[14967:14960] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[14975:14968] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[14983:14976] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[14991:14984] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[14999:14992] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[15007:15000] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[15015:15008] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[15023:15016] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[15031:15024] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[15039:15032] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[15047:15040] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[15055:15048] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[15063:15056] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[15071:15064] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[15079:15072] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[15087:15080] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[15095:15088] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[15103:15096] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[15111:15104] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[15119:15112] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[15127:15120] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[15135:15128] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[15143:15136] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[15151:15144] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[15159:15152] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[15167:15160] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[15175:15168] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[15183:15176] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[15191:15184] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[15199:15192] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[15207:15200] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[15215:15208] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[15223:15216] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[15231:15224] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[15239:15232] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[15247:15240] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[15255:15248] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[15263:15256] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[15271:15264] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[15279:15272] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[15287:15280] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[15295:15288] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[15303:15296] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[15311:15304] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[15319:15312] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[15327:15320] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[15335:15328] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[15343:15336] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[15351:15344] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[15359:15352] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[5].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[15367:15360] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[15375:15368] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[15383:15376] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[15391:15384] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[15399:15392] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[15407:15400] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[15415:15408] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[15423:15416] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[15431:15424] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[15439:15432] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[15447:15440] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[15455:15448] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[15463:15456] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[15471:15464] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[15479:15472] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[15487:15480] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[15495:15488] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[15503:15496] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[15511:15504] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[15519:15512] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[15527:15520] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[15535:15528] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[15543:15536] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[15551:15544] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[15559:15552] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[15567:15560] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[15575:15568] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[15583:15576] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[15591:15584] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[15599:15592] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[15607:15600] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[15615:15608] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[15623:15616] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[15631:15624] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[15639:15632] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[15647:15640] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[15655:15648] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[15663:15656] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[15671:15664] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[15679:15672] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[15687:15680] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[15695:15688] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[15703:15696] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[15711:15704] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[15719:15712] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[15727:15720] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[15735:15728] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[15743:15736] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[15751:15744] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[15759:15752] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[15767:15760] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[15775:15768] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[15783:15776] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[15791:15784] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[15799:15792] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[15807:15800] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[15815:15808] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[15823:15816] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[15831:15824] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[15839:15832] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[15847:15840] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[15855:15848] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[15863:15856] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[15871:15864] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[6].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[15879:15872] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[15887:15880] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[15895:15888] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[15903:15896] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[15911:15904] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[15919:15912] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[15927:15920] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[15935:15928] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[0].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[15943:15936] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[15951:15944] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[15959:15952] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[15967:15960] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[15975:15968] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[15983:15976] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[15991:15984] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[15999:15992] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[1].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[16007:16000] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[16015:16008] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[16023:16016] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[16031:16024] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[16039:16032] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[16047:16040] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[16055:16048] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[16063:16056] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[2].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[16071:16064] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[16079:16072] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[16087:16080] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[16095:16088] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[16103:16096] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[16111:16104] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[16119:16112] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[16127:16120] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[3].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[16135:16128] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[16143:16136] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[16151:16144] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[16159:16152] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[16167:16160] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[16175:16168] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[16183:16176] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[16191:16184] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[4].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[16199:16192] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[16207:16200] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[16215:16208] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[16223:16216] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[16231:16224] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[16239:16232] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[16247:16240] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[16255:16248] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[5].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[16263:16256] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[16271:16264] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[16279:16272] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[16287:16280] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[16295:16288] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[16303:16296] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[16311:16304] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[16319:16312] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[6].ram64_inst.genblk1[7].ram8_inst.mem;
 mem[16327:16320] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[0].ram8_inst.mem;
 mem[16335:16328] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[1].ram8_inst.mem;
 mem[16343:16336] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[2].ram8_inst.mem;
 mem[16351:16344] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[3].ram8_inst.mem;
 mem[16359:16352] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[4].ram8_inst.mem;
 mem[16367:16360] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[5].ram8_inst.mem;
 mem[16375:16368] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[6].ram8_inst.mem;
 mem[16383:16376] =dut.ram16k_inst.genblk1[3].ram4k_inst.genblk1[7].ram512_inst.genblk1[7].ram64_inst.genblk1[7].ram8_inst.mem;



end

 
// Stimulus
initial begin
// Initialize inputs

clk = 0;
reset = 0;

// Wait for a few clock cycles
#10;

// Deassert reset
reset = 1;

// write mem vector to file, to see what in memory
f1 = $fopen("tb_mem1.txt","w");
$fwrite(f1,"%h",mem);

// Wait for simulation to complete
#100000000;

$fwrite(f1,"%h",mem);
$fclose(f1);
$finish;

end


endmodule